module ui

import (
	glfw
)

pub fn start() {
	glfw.init_glfw()
}
