module layout

pub struct Menu {}
